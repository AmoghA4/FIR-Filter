`timescale 1ns/1ps

module ROM_SONG1(
    clk,
    address,
    data
    );
    
    parameter DATA_WIDTH = 8;
    parameter ADDR_WIDTH = 10;
    
    input clk;
    input [9:0] address;
    
    output reg signed [DATA_WIDTH-1:0] data;

    always @ (posedge clk)
    begin
        case(address)
            10'd0:   data <= 8'b00000000;
            10'd1:   data <= 8'b00000010;
            10'd2:   data <= 8'b00000100;
            10'd3:   data <= 8'b00000110;
            10'd4:   data <= 8'b00001000;
            10'd5:   data <= 8'b00001010;
            10'd6:   data <= 8'b00001100;
            10'd7:   data <= 8'b00001110;
            10'd8:   data <= 8'b00010000;
            10'd9:   data <= 8'b00010010;
            10'd10:  data <= 8'b00010010; 
            10'd11:  data <= 8'b00010100;
            10'd12:  data <= 8'b00010110;
            10'd13:  data <= 8'b00011000;
            10'd14:  data <= 8'b00011010;
            10'd15:  data <= 8'b00011100;
            10'd16:  data <= 8'b00011110;
            10'd17:  data <= 8'b00100000;
            10'd18:  data <= 8'b00100010;
            10'd19:  data <= 8'b00100011;            
            10'd20:  data <= 8'b00100101; 
            10'd21:  data <= 8'b00100111;
            10'd22:  data <= 8'b00101001;
            10'd23:  data <= 8'b00101011;
            10'd24:  data <= 8'b00101101;
            10'd25:  data <= 8'b00101111;            
            10'd26:  data <= 8'b00110001;
            10'd27:  data <= 8'b00110010;            
            10'd28:  data <= 8'b00110100;
            10'd29:  data <= 8'b00110110;            
            10'd30:  data <= 8'b00111000; 
            10'd31:  data <= 8'b00111010;
            10'd32:  data <= 8'b00111011;
            10'd33:  data <= 8'b00111101;
            10'd34:  data <= 8'b00111111;
            10'd35:  data <= 8'b01000001;            
            10'd36:  data <= 8'b01000010;
            10'd37:  data <= 8'b01000100;            
            10'd38:  data <= 8'b01000110;
            10'd39:  data <= 8'b01000111;
            
            10'd40:  data <= 8'b01001001; 
            10'd41:  data <= 8'b01001011;
            10'd42:  data <= 8'b01001100;
            10'd43:  data <= 8'b01001110;
            10'd44:  data <= 8'b01001111;
            10'd45:  data <= 8'b01010001;            
            10'd46:  data <= 8'b01010010;
            10'd47:  data <= 8'b01010100;            
            10'd48:  data <= 8'b01010101;
            10'd49:  data <= 8'b01010111;
            
            10'd50:  data <= 8'b01011000; 
            10'd51:  data <= 8'b01011010;
            10'd52:  data <= 8'b01011011;
            10'd53:  data <= 8'b01011101;
            10'd54:  data <= 8'b01011110;
            10'd55:  data <= 8'b01011111;            
            10'd56:  data <= 8'b01100001;
            10'd57:  data <= 8'b01100010;            
            10'd58:  data <= 8'b01100011;
            10'd59:  data <= 8'b01100100;
            
            10'd60:  data <= 8'b01100110; 
            10'd61:  data <= 8'b01100111;
            10'd62:  data <= 8'b01101000;
            10'd63:  data <= 8'b01101001;
            10'd64:  data <= 8'b01101010;
            10'd65:  data <= 8'b01101011;            
            10'd66:  data <= 8'b01101100;
            10'd67:  data <= 8'b01101101;            
            10'd68:  data <= 8'b01101110;
            10'd69:  data <= 8'b01101111;
            10'd70:  data <= 8'b01110000; 
            10'd71:  data <= 8'b01110001;
            10'd72:  data <= 8'b01110010;
            10'd73:  data <= 8'b01110011;            
            10'd74:  data <= 8'b01110100;
            10'd75:  data <= 8'b01110101;            
            10'd76:  data <= 8'b01110101;
            10'd77:  data <= 8'b01110110;            
            10'd78:  data <= 8'b01110111;
            10'd79:  data <= 8'b01110111;
            
            10'd80:  data <= 8'b01111000; 
            10'd81:  data <= 8'b01111001;
            10'd82:  data <= 8'b01111001;
            10'd83:  data <= 8'b01111010;
            10'd84:  data <= 8'b01111010;
            10'd85:  data <= 8'b01111011;            
            10'd86:  data <= 8'b01111011;
            10'd87:  data <= 8'b01111100;            
            10'd88:  data <= 8'b01111100;
            10'd89:  data <= 8'b01111101;        
            10'd90:  data <= 8'b01111101; 
            10'd91:  data <= 8'b01111101;
            10'd92:  data <= 8'b01111110;
            10'd93:  data <= 8'b01111110;
            10'd94:  data <= 8'b01111110;
            10'd95:  data <= 8'b01111110;            
            10'd96:  data <= 8'b01111111;
            10'd97:  data <= 8'b01111111;            
            10'd98:  data <= 8'b01111111;
            10'd99:  data <= 8'b01111111;            
            10'd100: data <= 8'b01111111; 
            10'd101: data <= 8'b01111111;
            10'd102: data <= 8'b01111111;
            10'd103: data <= 8'b01111111;
            10'd104: data <= 8'b01111111;
            10'd105: data <= 8'b01111111;            
            10'd106: data <= 8'b01111110;
            10'd107: data <= 8'b01111110;            
            10'd108: data <= 8'b01111110;
            10'd109: data <= 8'b01111110;            
            10'd110: data <= 8'b01111101; 
            10'd111: data <= 8'b01111101;
            10'd112: data <= 8'b01111101;
            10'd113: data <= 8'b01111100;
            10'd114: data <= 8'b01111100;
            10'd115: data <= 8'b01111011;            
            10'd116: data <= 8'b01111011;
            10'd117: data <= 8'b01111010;            
            10'd118: data <= 8'b01111010;
            10'd119: data <= 8'b01111001;            
            10'd120: data <= 8'b01111001; 
            10'd121: data <= 8'b01111000;
            10'd122: data <= 8'b01110111;
            10'd123: data <= 8'b01110111;
            10'd124: data <= 8'b01110110;
            10'd125: data <= 8'b01110101;            
            10'd126: data <= 8'b01110101;
            10'd127: data <= 8'b01110100;            
            10'd128: data <= 8'b01110011;
            10'd129: data <= 8'b01110010;            
            10'd130: data <= 8'b01110001; 
            10'd131: data <= 8'b01110000;
            10'd132: data <= 8'b01101111;
            10'd133: data <= 8'b01101110;
            10'd134: data <= 8'b01101101;
            10'd135: data <= 8'b01101100;            
            10'd136: data <= 8'b01101011;
            10'd137: data <= 8'b01101010;            
            10'd138: data <= 8'b01101001;
            10'd139: data <= 8'b01101000;            
            10'd140: data <= 8'b01100111; 
            10'd141: data <= 8'b01100110;
            10'd142: data <= 8'b01100100;
            10'd143: data <= 8'b01100011;
            10'd144: data <= 8'b01100010;
            10'd145: data <= 8'b01100001;            
            10'd146: data <= 8'b01011111;
            10'd147: data <= 8'b01011110;            
            10'd148: data <= 8'b01011101;
            10'd149: data <= 8'b01011011;            
            10'd150: data <= 8'b01011010; 
            10'd151: data <= 8'b01011000;
            10'd152: data <= 8'b01010111;
            10'd153: data <= 8'b01010101;
            10'd154: data <= 8'b01010100;
            10'd155: data <= 8'b01010010;            
            10'd156: data <= 8'b01010001;
            10'd157: data <= 8'b01001111;            
            10'd158: data <= 8'b01001110;
            10'd159: data <= 8'b01001100;
            
            10'd160: data <= 8'b01001011; 
            10'd161: data <= 8'b01001001;
            10'd162: data <= 8'b01000111;
            10'd163: data <= 8'b01000110;
            10'd164: data <= 8'b01000100;
            10'd165: data <= 8'b01000010;            
            10'd166: data <= 8'b01000001;
            10'd167: data <= 8'b00111111;            
            10'd168: data <= 8'b00111101;
            10'd169: data <= 8'b00111011;            
            10'd170: data <= 8'b00111010; 
            10'd171: data <= 8'b00111000;
            10'd172: data <= 8'b00110110;
            10'd173: data <= 8'b00110100;
            10'd174: data <= 8'b00110010;
            10'd175: data <= 8'b00110001;            
            10'd176: data <= 8'b00101111;
            10'd177: data <= 8'b00101101;            
            10'd178: data <= 8'b00101011;
            10'd179: data <= 8'b00101001;
        
            10'd180: data <= 8'b00100111; 
            10'd181: data <= 8'b00100101;
            10'd182: data <= 8'b00100011;
            10'd183: data <= 8'b00100010;
            10'd184: data <= 8'b00100000;
            10'd185: data <= 8'b00011110;            
            10'd186: data <= 8'b00011100;
            10'd187: data <= 8'b00011010;            
            10'd188: data <= 8'b00011000;
            10'd189: data <= 8'b00010110;

            10'd190: data <= 8'b00010100; 
            10'd191: data <= 8'b00010010;
            10'd192: data <= 8'b00010000;
            10'd193: data <= 8'b00001110;
            10'd194: data <= 8'b00001100;
            10'd195: data <= 8'b00001010;            
            10'd196: data <= 8'b00001000;
            10'd197: data <= 8'b00000110;            
            10'd198: data <= 8'b00000100;
            10'd199: data <= 8'b00000010;
            
            10'd200: data <= 8'b00000000;
            10'd201: data <= 8'b11111110; 
          10'd202: data <= 8'b11111100; 
          10'd203: data <= 8'b11111010; 
          10'd204: data <= 8'b11111000; 
          10'd205: data <= 8'b11110110; 
          10'd206: data <= 8'b11110100; 
          10'd207: data <= 8'b11110010; 
          10'd208: data <= 8'b11110000; 
          10'd209: data <= 8'b11101110; 
          10'd210: data <= 8'b11101100; 
          10'd211: data <= 8'b11101010; 
          10'd212: data <= 8'b11101000; 
          10'd213: data <= 8'b11100110; 
          10'd214: data <= 8'b11100100; 
          10'd215: data <= 8'b11100010;
          10'd216: data <= 8'b11100000;
          10'd217: data <= 8'b11011110;
          10'd218: data <= 8'b11011101;
          10'd219: data <= 8'b11011011;
          10'd220: data <= 8'b11011001;
          10'd221: data <= 8'b11010111;
          10'd222: data <= 8'b11010101;
          10'd223: data <= 8'b11010011;
          10'd224: data <= 8'b11010001;
          10'd225: data <= 8'b11001111;
          10'd226: data <= 8'b11001110;
          10'd227: data <= 8'b11001100;
          10'd228: data <= 8'b11001010;
          10'd229: data <= 8'b11001000;
          10'd230: data <= 8'b11000110;
          10'd231: data <= 8'b11000101;
          10'd232: data <= 8'b11000011;
          10'd233: data <= 8'b11000001;
          10'd234: data <= 8'b10111111;
          10'd235: data <= 8'b10111110; 
          10'd236: data <= 8'b10111100; 
          10'd237: data <= 8'b10111010; 
          10'd238: data <= 8'b10111001; 
          10'd239: data <= 8'b10110111; 
          10'd240: data <= 8'b10110101; 
          10'd241: data <= 8'b10110100; 
          10'd242: data <= 8'b10110010; 
          10'd243: data <= 8'b10110001; 
          10'd244: data <= 8'b10101111; 
          10'd245: data <= 8'b10101110; 
          10'd246: data <= 8'b10101110; 
          10'd247: data <= 8'b10101011; 
          10'd248: data <= 8'b10101001; 
          10'd249: data <= 8'b10101000; 
          10'd250: data <= 8'b10100110; 
          10'd251: data <= 8'b10100101; 
          10'd252: data <= 8'b10100011; 
          10'd253: data <= 8'b10100010; 
          10'd254: data <= 8'b10100001; 
          10'd255: data <= 8'b10011111; 
          10'd256: data <= 8'b10011110; 
          10'd257: data <= 8'b10011101; 
          10'd258: data <= 8'b10011100; 
          10'd259: data <= 8'b10011010; 
          10'd260: data <= 8'b10011001; 
          10'd261: data <= 8'b10011000; 
          10'd262: data <= 8'b10010111; 
          10'd263: data <= 8'b10010110; 
          10'd264: data <= 8'b10010101; 
          10'd265: data <= 8'b10010100; 
          10'd266: data <= 8'b10010011; 
          10'd267: data <= 8'b10010010; 
          10'd268: data <= 8'b10010001;
          10'd269: data <= 8'b10010000;
          10'd270: data <= 8'b10001111;
          10'd271: data <= 8'b10001110;
          10'd272: data <= 8'b10001101;
          10'd273: data <= 8'b10001100;
          10'd274: data <= 8'b10001011;
          10'd275: data <= 8'b10001011;
          10'd276: data <= 8'b10001010;
          10'd277: data <= 8'b10001001;
          10'd278: data <= 8'b10001001;
          10'd279: data <= 8'b10001000;
          10'd280: data <= 8'b10000111;
          10'd281: data <= 8'b10000111;
          10'd282: data <= 8'b10000110;
          10'd283: data <= 8'b10000101;
          10'd284: data <= 8'b10000101;
          10'd285: data <= 8'b10000101;
          10'd286: data <= 8'b10000100;
          10'd287: data <= 8'b10000100;
          10'd288: data <= 8'b10000011;
          10'd289: data <= 8'b10000011;
          10'd290: data <= 8'b10000011;
          10'd291: data <= 8'b10000010;
          10'd292: data <= 8'b10000010;
          10'd293: data <= 8'b10000010;
          10'd294: data <= 8'b10000010;
          10'd295: data <= 8'b10000001;
          10'd296: data <= 8'b10000001;
          10'd297: data <= 8'b10000001;
          10'd298: data <= 8'b10000001;
          10'd299: data <= 8'b10000001;
          10'd300: data <= 8'b10000001;
          10'd301: data <= 8'b10000001;
          10'd302: data <= 8'b10000001;
          10'd303: data <= 8'b10000001;
          10'd304: data <= 8'b10000001;
          10'd305: data <= 8'b10000001;
          10'd306: data <= 8'b10000010;
          10'd307: data <= 8'b10000010;
          10'd308: data <= 8'b10000010;
          10'd309: data <= 8'b10000010;
          10'd310: data <= 8'b10000011;
          10'd311: data <= 8'b10000011;
          10'd312: data <= 8'b10000011;
          10'd313: data <= 8'b10000100;
          10'd314: data <= 8'b10000100;
          10'd315: data <= 8'b10000101;
          10'd316: data <= 8'b10000101;
          10'd317: data <= 8'b10000101;
          10'd318: data <= 8'b10000110;
          10'd319: data <= 8'b10000111;
          10'd320: data <= 8'b10000111;
          10'd321: data <= 8'b10001000;
          10'd322: data <= 8'b10001001;
          10'd323: data <= 8'b10001001;
          10'd324: data <= 8'b10001010;
          10'd325: data <= 8'b10001011;
          10'd326: data <= 8'b10001011;
          10'd327: data <= 8'b10001100;
          10'd328: data <= 8'b10001101;
          10'd329: data <= 8'b10001110;
          10'd330: data <= 8'b10001111;
          10'd331: data <= 8'b10010000;
          10'd332: data <= 8'b10010001;
          10'd333: data <= 8'b10010010;
          10'd334: data <= 8'b10010011;
          10'd335: data <= 8'b10010100;
          10'd336: data <= 8'b10010101;
          10'd337: data <= 8'b10010110;
          10'd338: data <= 8'b10010111;
          10'd339: data <= 8'b10011000;
          10'd340: data <= 8'b10011001;
          10'd341: data <= 8'b10011010;
          10'd342: data <= 8'b10011100;
          10'd343: data <= 8'b10011101;
          10'd344: data <= 8'b10011110;
          10'd345: data <= 8'b10011111;
          10'd346: data <= 8'b10100001;
          10'd347: data <= 8'b10100010;
          10'd348: data <= 8'b10100011;
          10'd349: data <= 8'b10100101;
          10'd350: data <= 8'b10100110;
          10'd351: data <= 8'b10101000;
          10'd352: data <= 8'b10101001;
          10'd353: data <= 8'b10101011;
          10'd354: data <= 8'b10101100;
          10'd355: data <= 8'b10101110;
          10'd356: data <= 8'b10101111;
          10'd357: data <= 8'b10110001; 
          10'd358: data <= 8'b10110010; 
          10'd359: data <= 8'b10110100; 
          10'd360: data <= 8'b10110101; 
          10'd361: data <= 8'b10110111; 
          10'd362: data <= 8'b10111001; 
          10'd363: data <= 8'b10111010; 
          10'd364: data <= 8'b10111100; 
          10'd365: data <= 8'b10111110; 
          10'd366: data <= 8'b10111111; 
          10'd367: data <= 8'b11000001; 
          10'd368: data <= 8'b11000011; 
          10'd369: data <= 8'b11000101; 
          10'd370: data <= 8'b11000110; 
          10'd371: data <= 8'b11001000; 
          10'd372: data <= 8'b11001010; 
          10'd373: data <= 8'b11001100; 
          10'd374: data <= 8'b11001110; 
          10'd375: data <= 8'b11001111; 
          10'd376: data <= 8'b11010001; 
          10'd377: data <= 8'b11010011; 
          10'd378: data <= 8'b11010101; 
          10'd379: data <= 8'b11010111; 
          10'd380: data <= 8'b11011001; 
          10'd381: data <= 8'b11011011; 
          10'd382: data <= 8'b11011101; 
          10'd383: data <= 8'b11011110; 
          10'd384: data <= 8'b11100000; 
          10'd385: data <= 8'b11100010; 
          10'd386: data <= 8'b11100100; 
          10'd387: data <= 8'b11100110; 
          10'd388: data <= 8'b11101000; 
          10'd389: data <= 8'b11101010; 
          10'd390: data <= 8'b11101100; 
          10'd391: data <= 8'b11101110; 
          10'd392: data <= 8'b11110000; 
          10'd393: data <= 8'b11110010; 
          10'd394: data <= 8'b11110100; 
          10'd395: data <= 8'b11110110; 
          10'd396: data <= 8'b11111000; 
          10'd397: data <= 8'b11111010; 
          10'd398: data <= 8'b11111100; 
          10'd399: data <= 8'b11111110; 
          10'd400: data <= 8'b00000000;
          default: data <= 8'b00000000;
        endcase
    end
    
endmodule